--------------------------------------------------------------------------------
-- Company: 	Queen Mary University
-- Engineer: 	Michael Seltene : 120099030
-- 				Group : 7
-- Create Date:   14:48:24 10/14/2015
-- Design Name:   full_adder
-- Module Name:   full_adder_test_bench.vhd
-- Project Name:  Lab 1
-- Target Device: XCR3064xl-6pc44
-- Tool versions: Xilinx ISE	   7.104i and ModelSim XE III 6.0a starter 
-- Description:   full adder test bench
-- 
-- VHDL Test Bench Created by ISE for module: full_adder
-- 
-- Dependencies:  full_adder.vhd
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;
 
-- ENTITY
ENTITY full_adder_test_bench IS
END full_adder_test_bench;
 
-- ARCHITECTURE
ARCHITECTURE behavior OF full_adder_test_bench IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT full_adder
    PORT(
         a : IN  std_logic;
         b : IN  std_logic;
         cin : IN  std_logic;
         s : OUT  std_logic;
         cout : OUT  std_logic
        );
    END COMPONENT;
    
   --Inputs
   signal a : std_logic := '0';
   signal b : std_logic := '0';
   signal cin : std_logic := '0';

 	--Outputs
   signal s : std_logic;
   signal cout : std_logic;
  
BEGIN
	-- Instantiate the Unit Under Test (UUT)
   uut: full_adder PORT MAP (
          a => a,
          b => b,
          cin => cin,
          s => s,
          cout => cout
        );


	   -- TRUTH TABLE --
-- ********************** --

--  a  b  cin  : s  cout
---------------:--------
--  0	 0	 0    : 0  0
--	 0	 0	 1    : 0  1
--	 0	 1	 0    : 0  1
--	 0	 1	 1    : 1  0
--	 1	 0	 0    : 0  1
--	 1	 0	 1    : 1  0
--	 1	 1	 0    : 1  0
--	 1	 1	 1    : 1  1

-- ********************** --

   -- Stimulus process
   stim_proc: process
   begin		
      -- Wait 100 ns for global reset to finish
		wait for 100 ns;
		a <= '0'; b <= '0'; cin <= '0'; 		-- check that 0 + 0 + 0 => cout = 0 sum = 0 	
		wait for 100 ns;
		a <= '1'; b <= '0'; cin <= '0'; 		-- check that 1 + 0 + 0 => cout = 0 sum = 1 	
		wait for 100 ns;
		a <= '0'; b <= '1'; cin <= '0'; 		-- check that 1 + 0 + 0 => cout = 0 sum = 1 	
		wait for 100 ns;
		a <= '1'; b <= '1'; cin <= '0'; 		-- check that 1 + 1 + 0 => cout = 1 sum = 0		
	   wait for 100 ns;
		a <= '0'; b <= '0'; cin <= '1'; 		-- check that 0 + 0 + 1 => cout = 0 sum = 1
		wait for 100 ns;
		a <= '1'; b <= '0'; cin <= '1'; 		-- check that 1 + 0 +  1 => cout = 1 sum = 0
		wait for 100 ns;
		a <= '0'; b <= '1'; cin <= '1'; 		-- check that 0 + 1 +  1 => cout = 1 sum = 0
		wait for 100 ns;
		a <= '1'; b <= '1'; cin <= '1'; 		-- check that 1 + 1 +  1 => cout = 1 sum = 1 
 
		wait; -- will wait forever
   end process;

END;
