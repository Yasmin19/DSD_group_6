----------------------------------------------------------------------------------
-- Company: 	QMUL
-- Engineer: 	Michael Seltene
-- 
-- Create Date:    12:55:57 11/24/2015 
-- Design Name: 	 tdm_display_circuit
-- Module Name:    tdm_display_circuit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity tdm_display_circuit is
end tdm_display_circuit;

architecture Behavioral of tdm_display_circuit is
	
begin


end Behavioral;

